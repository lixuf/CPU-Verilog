`timescale 1ns/1ps

module testbench;







reg [31:0] r_in;//输入指令

initial begin
r_in<=32'b01000100110001111101100100010110;
#5
r_in<=32'b01000011010000100010100110001010;
#5
r_in<=32'b00111111011001010011001100100010;
#5
r_in<=32'b01010110110010000111110100110011;
#5
r_in<=32'b00111011011111010011011011111101;
#5
r_in<=32'b00111101010111100100110111110011;
#5
r_in<=32'b01011000001100000011010110111001;
#5
r_in<=32'b00111001101111001110111101111111;
#5
r_in<=32'b00000001101010101010011101011100;
#5
r_in<=32'b00000011001001010100010101101011;
#5
r_in<=32'b00000100111010101010110000010101;
#5
r_in<=32'b00000110111100010101111001110111;
#5
r_in<=32'b00001000010101001000001000010101;
#5
r_in<=32'b00001010101111100100000101101111;
#5
r_in<=32'b00001100101110000000011100100111;
#5
r_in<=32'b00001110010111001001101001000010;
#5
r_in<=32'b00010001010000010111010101110010;
#5
r_in<=32'b00010010000101100100110111110110;
#5
r_in<=32'b00010100100010110010001000100011;
#5
r_in<=32'b00010110101111101011011111100100;
#5
r_in<=32'b00011000100001101100011010000000;
#5
r_in<=32'b00011010011100100101110101010010;
#5
r_in<=32'b00011101000000100000010010110100;
#5
r_in<=32'b00011110010001100001111011100100;
#5
r_in<=32'b00100001110100011000010100000101;
#5
r_in<=32'b00100011110001011100011111010001;
#5
r_in<=32'b00100100101000011101110100111000;
#5
r_in<=32'b00100111100101001010101101010101;
#5
r_in<=32'b00101001111010001110011000111011;
#5
r_in<=32'b00101010011001000010111100001110;
#5
r_in<=32'b00101100010000000101100000111000;
#5
r_in<=32'b00101111101110110101100001010000;
#5
r_in<=32'b00110001100100000101111110011101;
#5
r_in<=32'b00110010101111010001101110100000;
#5
r_in<=32'b00110101100001010011010010000100;
#5
r_in<=32'b00110111110000111001100111001100;
#5
r_in<=32'b01000001110111010110111111101000;
#5
r_in<=32'b01000110101011011001111010101001;
#5
r_in<=32'b01001000101101111000110110000001;
#5
r_in<=32'b01001010101101100100001100001110;
#5
r_in<=32'b01001100110011101111110101101001;
#5
r_in<=32'b01001110010101110101101010000101;
#5
r_in<=32'b01010001011000001101011110101011;
#5
r_in<=32'b01010010010110111111001100001110;
#5
r_in<=32'b01010101111001010111100101101110;
$stop;
end

//输出的控制信号
//修改寄存器
wire [7:0] xbh_en;//在一级流水处锁存
wire [7:0] xbl_en;
wire [7:0] fir_reg_en;
wire [1:0] des_addr_en;
wire [1:0] sor_addr_en;
wire len_en;
wire [3:0] lr_en;
wire [3:0] hr_en;
wire [15:0] operand;
//指令部分
////ad
wire ad_en;
wire des;
wire [7:0] select;
////小波分解;fir滤波器指令;uart输出指令
wire xb_en;
wire fir_en;
wire uarto_en;
wire [7:0] channel;//控制ad通道
wire [1:0] source;//介质选择 10 ad 00 ram 01 ddr
//wire [7:0] select;
////中值滤波指令
wire zlb_en;
//wire [1:0] source;
////存储器搬移指令
wire move_en;
wire dir;
////中断等待指令
wire int_en;
////检测器启用指令
wire jc_en;
//wire [7:0] channel,



decoder dec(
.r_in(r_in),//输入指令


//输出的控制信号
//修改寄存器
.xbh_en(xbh_en),//在一级流水处锁存
.xbl_en(xbl_en),
. fir_reg_en(fir_reg_en),
. des_addr_en(des_addr_en),
. sor_addr_en(sor_addr_en),
. len_en(len_en),
. lr_en(lr_en),
. hr_en(hr_en),
.  operand(operand),
//指令部分
////ad
. ad_en(ad_en),
. des(des),
.  select(select),
////小波分解,fir滤波器指令,uart输出指令
. xb_en(xb_en),
. fir_en(fir_en),
. uarto_en(uarto_en),
. channel(channel),//控制ad通道
. source(source),//介质选择 10 ad 00 ram 01 ddr
//. [7:0] select,
////中值滤波指令
. zlb_en(zlb_en),
//. [1:0] source,
////存储器搬移指令
. move_en(move_en),
. dir(dir),
////中断等待指令
. int_en( int_en),
////检测( int_en器启用指令
. jc_en(jc_en)
//. [7:0] channel,


);







endmodule
